module Font_ROM(
  input logic clk,
  input logic [11:0] address, //Pendiente: Agregar ASCII extendido
  output logic [7:0] data
);
  logic [7:0] font [0:2019];

  always @ (posedge clk) begin
    if (address > 11'h7e3)
      data <= 8'h0;
    else
      data <= font[address];
  end

  initial begin
    font[0] = 8'h0;
    font[1] = 8'h0;
    font[2] = 8'h66;
    font[3] = 8'h42;
    font[4] = 8'h0;
    font[5] = 8'h42;
    font[6] = 8'h42;
    font[7] = 8'h42;
    font[8] = 8'h0;
    font[9] = 8'h42;
    font[10] = 8'h42;
    font[11] = 8'h66;
    font[12] = 8'h0;
    font[13] = 8'h0;
    font[14] = 8'h0;
    font[15] = 8'h0;
    font[16] = 8'h0;
    font[17] = 8'h0;
    font[18] = 8'h0;
    font[19] = 8'h0;
    font[20] = 8'h0;
    font[21] = 8'h0;
    font[22] = 8'h0;
    font[23] = 8'h0;
    font[24] = 8'h0;
    font[25] = 8'h0;
    font[26] = 8'h0;
    font[27] = 8'h0;
    font[28] = 8'h0;
    font[29] = 8'h0;
    font[30] = 8'h0;
    font[31] = 8'h0;
    font[32] = 8'h0;
    font[33] = 8'h0;
    font[34] = 8'h0;
    font[35] = 8'h0;
    font[36] = 8'h0;
    font[37] = 8'h0;
    font[38] = 8'h0;
    font[39] = 8'h0;
    font[40] = 8'h0;
    font[41] = 8'h0;
    font[42] = 8'h0;
    font[43] = 8'h0;
    font[44] = 8'h0;
    font[45] = 8'h0;
    font[46] = 8'h0;
    font[47] = 8'h0;
    font[48] = 8'h0;
    font[49] = 8'h0;
    font[50] = 8'h0;
    font[51] = 8'h0;
    font[52] = 8'h0;
    font[53] = 8'h0;
    font[54] = 8'h0;
    font[55] = 8'h0;
    font[56] = 8'h0;
    font[57] = 8'h0;
    font[58] = 8'h0;
    font[59] = 8'h0;
    font[60] = 8'h0;
    font[61] = 8'h0;
    font[62] = 8'h0;
    font[63] = 8'h0;
    font[64] = 8'h0;
    font[65] = 8'h0;
    font[66] = 8'h0;
    font[67] = 8'h0;
    font[68] = 8'h0;
    font[69] = 8'h0;
    font[70] = 8'h0;
    font[71] = 8'h0;
    font[72] = 8'h0;
    font[73] = 8'h0;
    font[74] = 8'h0;
    font[75] = 8'h0;
    font[76] = 8'h0;
    font[77] = 8'h0;
    font[78] = 8'h0;
    font[79] = 8'h0;
    font[80] = 8'h0;
    font[81] = 8'h0;
    font[82] = 8'h0;
    font[83] = 8'h0;
    font[84] = 8'h0;
    font[85] = 8'h0;
    font[86] = 8'h0;
    font[87] = 8'h0;
    font[88] = 8'h0;
    font[89] = 8'h0;
    font[90] = 8'h0;
    font[91] = 8'h0;
    font[92] = 8'h0;
    font[93] = 8'h0;
    font[94] = 8'h0;
    font[95] = 8'h0;
    font[96] = 8'h0;
    font[97] = 8'h0;
    font[98] = 8'h0;
    font[99] = 8'h0;
    font[100] = 8'h0;
    font[101] = 8'h0;
    font[102] = 8'h0;
    font[103] = 8'h0;
    font[104] = 8'h0;
    font[105] = 8'h0;
    font[106] = 8'h0;
    font[107] = 8'h0;
    font[108] = 8'h0;
    font[109] = 8'h0;
    font[110] = 8'h0;
    font[111] = 8'h0;
    font[112] = 8'h0;
    font[113] = 8'h0;
    font[114] = 8'h0;
    font[115] = 8'h0;
    font[116] = 8'h0;
    font[117] = 8'h0;
    font[118] = 8'h0;
    font[119] = 8'h0;
    font[120] = 8'h0;
    font[121] = 8'h0;
    font[122] = 8'h0;
    font[123] = 8'h0;
    font[124] = 8'h0;
    font[125] = 8'h0;
    font[126] = 8'h0;
    font[127] = 8'h0;
    font[128] = 8'h0;
    font[129] = 8'h0;
    font[130] = 8'h0;
    font[131] = 8'h0;
    font[132] = 8'h0;
    font[133] = 8'h0;
    font[134] = 8'h0;
    font[135] = 8'h0;
    font[136] = 8'h0;
    font[137] = 8'h0;
    font[138] = 8'h0;
    font[139] = 8'h0;
    font[140] = 8'h0;
    font[141] = 8'h0;
    font[142] = 8'h0;
    font[143] = 8'h0;
    font[144] = 8'h0;
    font[145] = 8'h0;
    font[146] = 8'h0;
    font[147] = 8'h0;
    font[148] = 8'h0;
    font[149] = 8'h0;
    font[150] = 8'h0;
    font[151] = 8'h0;
    font[152] = 8'h0;
    font[153] = 8'h0;
    font[154] = 8'h0;
    font[155] = 8'h0;
    font[156] = 8'h0;
    font[157] = 8'h0;
    font[158] = 8'h0;
    font[159] = 8'h0;
    font[160] = 8'h0;
    font[161] = 8'h0;
    font[162] = 8'h0;
    font[163] = 8'h0;
    font[164] = 8'h0;
    font[165] = 8'h0;
    font[166] = 8'h0;
    font[167] = 8'h0;
    font[168] = 8'h0;
    font[169] = 8'h0;
    font[170] = 8'h0;
    font[171] = 8'h0;
    font[172] = 8'h0;
    font[173] = 8'h0;
    font[174] = 8'h0;
    font[175] = 8'h0;
    font[176] = 8'h0;
    font[177] = 8'h0;
    font[178] = 8'h0;
    font[179] = 8'h0;
    font[180] = 8'h0;
    font[181] = 8'h0;
    font[182] = 8'h0;
    font[183] = 8'h0;
    font[184] = 8'h0;
    font[185] = 8'h0;
    font[186] = 8'h0;
    font[187] = 8'h0;
    font[188] = 8'h0;
    font[189] = 8'h0;
    font[190] = 8'h0;
    font[191] = 8'h0;
    font[192] = 8'h0;
    font[193] = 8'h0;
    font[194] = 8'h0;
    font[195] = 8'h0;
    font[196] = 8'h0;
    font[197] = 8'h0;
    font[198] = 8'h0;
    font[199] = 8'h0;
    font[200] = 8'h0;
    font[201] = 8'h0;
    font[202] = 8'h0;
    font[203] = 8'h0;
    font[204] = 8'h0;
    font[205] = 8'h0;
    font[206] = 8'h0;
    font[207] = 8'h0;
    font[208] = 8'h0;
    font[209] = 8'h0;
    font[210] = 8'h0;
    font[211] = 8'h0;
    font[212] = 8'h0;
    font[213] = 8'h0;
    font[214] = 8'h0;
    font[215] = 8'h0;
    font[216] = 8'h0;
    font[217] = 8'h0;
    font[218] = 8'h0;
    font[219] = 8'h0;
    font[220] = 8'h0;
    font[221] = 8'h0;
    font[222] = 8'h0;
    font[223] = 8'h0;
    font[224] = 8'h0;
    font[225] = 8'h0;
    font[226] = 8'h0;
    font[227] = 8'h0;
    font[228] = 8'h0;
    font[229] = 8'h0;
    font[230] = 8'h0;
    font[231] = 8'h0;
    font[232] = 8'h0;
    font[233] = 8'h0;
    font[234] = 8'h0;
    font[235] = 8'h0;
    font[236] = 8'h0;
    font[237] = 8'h0;
    font[238] = 8'h0;
    font[239] = 8'h0;
    font[240] = 8'h0;
    font[241] = 8'h0;
    font[242] = 8'h0;
    font[243] = 8'h0;
    font[244] = 8'h0;
    font[245] = 8'h0;
    font[246] = 8'h0;
    font[247] = 8'h0;
    font[248] = 8'h0;
    font[249] = 8'h0;
    font[250] = 8'h0;
    font[251] = 8'h0;
    font[252] = 8'h0;
    font[253] = 8'h0;
    font[254] = 8'h0;
    font[255] = 8'h0;
    font[256] = 8'h0;
    font[257] = 8'h0;
    font[258] = 8'h0;
    font[259] = 8'h0;
    font[260] = 8'h0;
    font[261] = 8'h0;
    font[262] = 8'h0;
    font[263] = 8'h0;
    font[264] = 8'h0;
    font[265] = 8'h0;
    font[266] = 8'h0;
    font[267] = 8'h0;
    font[268] = 8'h0;
    font[269] = 8'h0;
    font[270] = 8'h0;
    font[271] = 8'h0;
    font[272] = 8'h0;
    font[273] = 8'h0;
    font[274] = 8'h0;
    font[275] = 8'h0;
    font[276] = 8'h0;
    font[277] = 8'h0;
    font[278] = 8'h0;
    font[279] = 8'h0;
    font[280] = 8'h0;
    font[281] = 8'h0;
    font[282] = 8'h0;
    font[283] = 8'h0;
    font[284] = 8'h0;
    font[285] = 8'h0;
    font[286] = 8'h0;
    font[287] = 8'h0;
    font[288] = 8'h0;
    font[289] = 8'h0;
    font[290] = 8'h0;
    font[291] = 8'h0;
    font[292] = 8'h0;
    font[293] = 8'h0;
    font[294] = 8'h0;
    font[295] = 8'h0;
    font[296] = 8'h0;
    font[297] = 8'h0;
    font[298] = 8'h0;
    font[299] = 8'h0;
    font[300] = 8'h0;
    font[301] = 8'h0;
    font[302] = 8'h0;
    font[303] = 8'h0;
    font[304] = 8'h0;
    font[305] = 8'h0;
    font[306] = 8'h0;
    font[307] = 8'h0;
    font[308] = 8'h0;
    font[309] = 8'h0;
    font[310] = 8'h0;
    font[311] = 8'h0;
    font[312] = 8'h0;
    font[313] = 8'h0;
    font[314] = 8'h0;
    font[315] = 8'h0;
    font[316] = 8'h0;
    font[317] = 8'h0;
    font[318] = 8'h0;
    font[319] = 8'h0;
    font[320] = 8'h0;
    font[321] = 8'h0;
    font[322] = 8'h0;
    font[323] = 8'h0;
    font[324] = 8'h0;
    font[325] = 8'h0;
    font[326] = 8'h0;
    font[327] = 8'h0;
    font[328] = 8'h0;
    font[329] = 8'h0;
    font[330] = 8'h0;
    font[331] = 8'h0;
    font[332] = 8'h0;
    font[333] = 8'h0;
    font[334] = 8'h0;
    font[335] = 8'h0;
    font[336] = 8'h0;
    font[337] = 8'h0;
    font[338] = 8'h0;
    font[339] = 8'h0;
    font[340] = 8'h0;
    font[341] = 8'h0;
    font[342] = 8'h0;
    font[343] = 8'h0;
    font[344] = 8'h0;
    font[345] = 8'h0;
    font[346] = 8'h0;
    font[347] = 8'h0;
    font[348] = 8'h0;
    font[349] = 8'h0;
    font[350] = 8'h0;
    font[351] = 8'h0;
    font[352] = 8'h0;
    font[353] = 8'h0;
    font[354] = 8'h0;
    font[355] = 8'h0;
    font[356] = 8'h0;
    font[357] = 8'h0;
    font[358] = 8'h0;
    font[359] = 8'h0;
    font[360] = 8'h0;
    font[361] = 8'h0;
    font[362] = 8'h0;
    font[363] = 8'h0;
    font[364] = 8'h0;
    font[365] = 8'h0;
    font[366] = 8'h0;
    font[367] = 8'h0;
    font[368] = 8'h0;
    font[369] = 8'h0;
    font[370] = 8'h0;
    font[371] = 8'h0;
    font[372] = 8'h0;
    font[373] = 8'h0;
    font[374] = 8'h0;
    font[375] = 8'h0;
    font[376] = 8'h0;
    font[377] = 8'h0;
    font[378] = 8'h0;
    font[379] = 8'h0;
    font[380] = 8'h0;
    font[381] = 8'h0;
    font[382] = 8'h0;
    font[383] = 8'h0;
    font[384] = 8'h0;
    font[385] = 8'h0;
    font[386] = 8'h0;
    font[387] = 8'h0;
    font[388] = 8'h0;
    font[389] = 8'h0;
    font[390] = 8'h0;
    font[391] = 8'h0;
    font[392] = 8'h0;
    font[393] = 8'h0;
    font[394] = 8'h0;
    font[395] = 8'h0;
    font[396] = 8'h0;
    font[397] = 8'h0;
    font[398] = 8'h0;
    font[399] = 8'h0;
    font[400] = 8'h0;
    font[401] = 8'h0;
    font[402] = 8'h0;
    font[403] = 8'h0;
    font[404] = 8'h0;
    font[405] = 8'h0;
    font[406] = 8'h0;
    font[407] = 8'h0;
    font[408] = 8'h0;
    font[409] = 8'h0;
    font[410] = 8'h0;
    font[411] = 8'h0;
    font[412] = 8'h0;
    font[413] = 8'h0;
    font[414] = 8'h0;
    font[415] = 8'h0;
    font[416] = 8'h0;
    font[417] = 8'h0;
    font[418] = 8'h0;
    font[419] = 8'h0;
    font[420] = 8'h0;
    font[421] = 8'h0;
    font[422] = 8'h0;
    font[423] = 8'h0;
    font[424] = 8'h0;
    font[425] = 8'h0;
    font[426] = 8'h0;
    font[427] = 8'h0;
    font[428] = 8'h0;
    font[429] = 8'h0;
    font[430] = 8'h0;
    font[431] = 8'h0;
    font[432] = 8'h0;
    font[433] = 8'h0;
    font[434] = 8'h0;
    font[435] = 8'h0;
    font[436] = 8'h0;
    font[437] = 8'h0;
    font[438] = 8'h0;
    font[439] = 8'h0;
    font[440] = 8'h0;
    font[441] = 8'h0;
    font[442] = 8'h0;
    font[443] = 8'h0;
    font[444] = 8'h0;
    font[445] = 8'h0;
    font[446] = 8'h0;
    font[447] = 8'h0;
    font[448] = 8'h0;
    font[449] = 8'h0;
    font[450] = 8'h0;
    font[451] = 8'h0;
    font[452] = 8'h0;
    font[453] = 8'h0;
    font[454] = 8'h0;
    font[455] = 8'h0;
    font[456] = 8'h0;
    font[457] = 8'h0;
    font[458] = 8'h0;
    font[459] = 8'h0;
    font[460] = 8'h0;
    font[461] = 8'h0;
    font[462] = 8'h0;
    font[463] = 8'h0;
    font[464] = 8'h0;
    font[465] = 8'h0;
    font[466] = 8'h0;
    font[467] = 8'h0;
    font[468] = 8'h0;
    font[469] = 8'h0;
    font[470] = 8'h0;
    font[471] = 8'h0;
    font[472] = 8'h0;
    font[473] = 8'h0;
    font[474] = 8'h0;
    font[475] = 8'h0;
    font[476] = 8'h0;
    font[477] = 8'h0;
    font[478] = 8'h0;
    font[479] = 8'h0;
    font[480] = 8'h0;
    font[481] = 8'h0;
    font[482] = 8'h0;
    font[483] = 8'h0;
    font[484] = 8'h0;
    font[485] = 8'h0;
    font[486] = 8'h0;
    font[487] = 8'h0;
    font[488] = 8'h0;
    font[489] = 8'h0;
    font[490] = 8'h0;
    font[491] = 8'h0;
    font[492] = 8'h0;
    font[493] = 8'h0;
    font[494] = 8'h0;
    font[495] = 8'h0;
    font[496] = 8'h0;
    font[497] = 8'h0;
    font[498] = 8'h0;
    font[499] = 8'h0;
    font[500] = 8'h0;
    font[501] = 8'h0;
    font[502] = 8'h0;
    font[503] = 8'h0;
    font[504] = 8'h0;
    font[505] = 8'h0;
    font[506] = 8'h0;
    font[507] = 8'h0;
    font[508] = 8'h0;
    font[509] = 8'h0;
    font[510] = 8'h0;
    font[511] = 8'h0;
    font[512] = 8'h0;
    font[513] = 8'h0;
    font[514] = 8'h0;
    font[515] = 8'h0;
    font[516] = 8'h0;
    font[517] = 8'h0;
    font[518] = 8'h0;
    font[519] = 8'h0;
    font[520] = 8'h0;
    font[521] = 8'h0;
    font[522] = 8'h0;
    font[523] = 8'h0;
    font[524] = 8'h0;
    font[525] = 8'h0;
    font[526] = 8'h0;
    font[527] = 8'h0;
    font[528] = 8'h0;
    font[529] = 8'h0;
    font[530] = 8'h10;
    font[531] = 8'h10;
    font[532] = 8'h10;
    font[533] = 8'h10;
    font[534] = 8'h10;
    font[535] = 8'h10;
    font[536] = 8'h10;
    font[537] = 8'h0;
    font[538] = 8'h10;
    font[539] = 8'h10;
    font[540] = 8'h0;
    font[541] = 8'h0;
    font[542] = 8'h0;
    font[543] = 8'h0;
    font[544] = 8'h0;
    font[545] = 8'h24;
    font[546] = 8'h24;
    font[547] = 8'h24;
    font[548] = 8'h0;
    font[549] = 8'h0;
    font[550] = 8'h0;
    font[551] = 8'h0;
    font[552] = 8'h0;
    font[553] = 8'h0;
    font[554] = 8'h0;
    font[555] = 8'h0;
    font[556] = 8'h0;
    font[557] = 8'h0;
    font[558] = 8'h0;
    font[559] = 8'h0;
    font[560] = 8'h0;
    font[561] = 8'h0;
    font[562] = 8'h24;
    font[563] = 8'h24;
    font[564] = 8'h24;
    font[565] = 8'h7e;
    font[566] = 8'h24;
    font[567] = 8'h24;
    font[568] = 8'h7e;
    font[569] = 8'h24;
    font[570] = 8'h24;
    font[571] = 8'h24;
    font[572] = 8'h0;
    font[573] = 8'h0;
    font[574] = 8'h0;
    font[575] = 8'h0;
    font[576] = 8'h0;
    font[577] = 8'h10;
    font[578] = 8'h10;
    font[579] = 8'h7c;
    font[580] = 8'h92;
    font[581] = 8'h90;
    font[582] = 8'h90;
    font[583] = 8'h7c;
    font[584] = 8'h12;
    font[585] = 8'h12;
    font[586] = 8'h92;
    font[587] = 8'h7c;
    font[588] = 8'h10;
    font[589] = 8'h10;
    font[590] = 8'h0;
    font[591] = 8'h0;
    font[592] = 8'h0;
    font[593] = 8'h0;
    font[594] = 8'h64;
    font[595] = 8'h94;
    font[596] = 8'h68;
    font[597] = 8'h8;
    font[598] = 8'h10;
    font[599] = 8'h10;
    font[600] = 8'h20;
    font[601] = 8'h2c;
    font[602] = 8'h52;
    font[603] = 8'h4c;
    font[604] = 8'h0;
    font[605] = 8'h0;
    font[606] = 8'h0;
    font[607] = 8'h0;
    font[608] = 8'h0;
    font[609] = 8'h0;
    font[610] = 8'h18;
    font[611] = 8'h24;
    font[612] = 8'h24;
    font[613] = 8'h18;
    font[614] = 8'h30;
    font[615] = 8'h4a;
    font[616] = 8'h44;
    font[617] = 8'h44;
    font[618] = 8'h44;
    font[619] = 8'h3a;
    font[620] = 8'h0;
    font[621] = 8'h0;
    font[622] = 8'h0;
    font[623] = 8'h0;
    font[624] = 8'h0;
    font[625] = 8'h10;
    font[626] = 8'h10;
    font[627] = 8'h10;
    font[628] = 8'h0;
    font[629] = 8'h0;
    font[630] = 8'h0;
    font[631] = 8'h0;
    font[632] = 8'h0;
    font[633] = 8'h0;
    font[634] = 8'h0;
    font[635] = 8'h0;
    font[636] = 8'h0;
    font[637] = 8'h0;
    font[638] = 8'h0;
    font[639] = 8'h0;
    font[640] = 8'h0;
    font[641] = 8'h0;
    font[642] = 8'h8;
    font[643] = 8'h10;
    font[644] = 8'h20;
    font[645] = 8'h20;
    font[646] = 8'h20;
    font[647] = 8'h20;
    font[648] = 8'h20;
    font[649] = 8'h20;
    font[650] = 8'h10;
    font[651] = 8'h8;
    font[652] = 8'h0;
    font[653] = 8'h0;
    font[654] = 8'h0;
    font[655] = 8'h0;
    font[656] = 8'h0;
    font[657] = 8'h0;
    font[658] = 8'h20;
    font[659] = 8'h10;
    font[660] = 8'h8;
    font[661] = 8'h8;
    font[662] = 8'h8;
    font[663] = 8'h8;
    font[664] = 8'h8;
    font[665] = 8'h8;
    font[666] = 8'h10;
    font[667] = 8'h20;
    font[668] = 8'h0;
    font[669] = 8'h0;
    font[670] = 8'h0;
    font[671] = 8'h0;
    font[672] = 8'h0;
    font[673] = 8'h0;
    font[674] = 8'h0;
    font[675] = 8'h0;
    font[676] = 8'h0;
    font[677] = 8'h24;
    font[678] = 8'h18;
    font[679] = 8'h7e;
    font[680] = 8'h18;
    font[681] = 8'h24;
    font[682] = 8'h0;
    font[683] = 8'h0;
    font[684] = 8'h0;
    font[685] = 8'h0;
    font[686] = 8'h0;
    font[687] = 8'h0;
    font[688] = 8'h0;
    font[689] = 8'h0;
    font[690] = 8'h0;
    font[691] = 8'h0;
    font[692] = 8'h0;
    font[693] = 8'h10;
    font[694] = 8'h10;
    font[695] = 8'h7c;
    font[696] = 8'h10;
    font[697] = 8'h10;
    font[698] = 8'h0;
    font[699] = 8'h0;
    font[700] = 8'h0;
    font[701] = 8'h0;
    font[702] = 8'h0;
    font[703] = 8'h0;
    font[704] = 8'h0;
    font[705] = 8'h0;
    font[706] = 8'h0;
    font[707] = 8'h0;
    font[708] = 8'h0;
    font[709] = 8'h0;
    font[710] = 8'h0;
    font[711] = 8'h0;
    font[712] = 8'h0;
    font[713] = 8'h0;
    font[714] = 8'h10;
    font[715] = 8'h10;
    font[716] = 8'h20;
    font[717] = 8'h0;
    font[718] = 8'h0;
    font[719] = 8'h0;
    font[720] = 8'h0;
    font[721] = 8'h0;
    font[722] = 8'h0;
    font[723] = 8'h0;
    font[724] = 8'h0;
    font[725] = 8'h0;
    font[726] = 8'h0;
    font[727] = 8'h7e;
    font[728] = 8'h0;
    font[729] = 8'h0;
    font[730] = 8'h0;
    font[731] = 8'h0;
    font[732] = 8'h0;
    font[733] = 8'h0;
    font[734] = 8'h0;
    font[735] = 8'h0;
    font[736] = 8'h0;
    font[737] = 8'h0;
    font[738] = 8'h0;
    font[739] = 8'h0;
    font[740] = 8'h0;
    font[741] = 8'h0;
    font[742] = 8'h0;
    font[743] = 8'h0;
    font[744] = 8'h0;
    font[745] = 8'h0;
    font[746] = 8'h10;
    font[747] = 8'h10;
    font[748] = 8'h0;
    font[749] = 8'h0;
    font[750] = 8'h0;
    font[751] = 8'h0;
    font[752] = 8'h0;
    font[753] = 8'h0;
    font[754] = 8'h4;
    font[755] = 8'h4;
    font[756] = 8'h8;
    font[757] = 8'h8;
    font[758] = 8'h10;
    font[759] = 8'h10;
    font[760] = 8'h20;
    font[761] = 8'h20;
    font[762] = 8'h40;
    font[763] = 8'h40;
    font[764] = 8'h0;
    font[765] = 8'h0;
    font[766] = 8'h0;
    font[767] = 8'h0;
    font[768] = 8'h0;
    font[769] = 8'h0;
    font[770] = 8'h3c;
    font[771] = 8'h42;
    font[772] = 8'h42;
    font[773] = 8'h46;
    font[774] = 8'h4a;
    font[775] = 8'h52;
    font[776] = 8'h62;
    font[777] = 8'h42;
    font[778] = 8'h42;
    font[779] = 8'h3c;
    font[780] = 8'h0;
    font[781] = 8'h0;
    font[782] = 8'h0;
    font[783] = 8'h0;
    font[784] = 8'h0;
    font[785] = 8'h0;
    font[786] = 8'h8;
    font[787] = 8'h18;
    font[788] = 8'h28;
    font[789] = 8'h8;
    font[790] = 8'h8;
    font[791] = 8'h8;
    font[792] = 8'h8;
    font[793] = 8'h8;
    font[794] = 8'h8;
    font[795] = 8'h3e;
    font[796] = 8'h0;
    font[797] = 8'h0;
    font[798] = 8'h0;
    font[799] = 8'h0;
    font[800] = 8'h0;
    font[801] = 8'h0;
    font[802] = 8'h3c;
    font[803] = 8'h42;
    font[804] = 8'h42;
    font[805] = 8'h2;
    font[806] = 8'h4;
    font[807] = 8'h8;
    font[808] = 8'h10;
    font[809] = 8'h20;
    font[810] = 8'h40;
    font[811] = 8'h7e;
    font[812] = 8'h0;
    font[813] = 8'h0;
    font[814] = 8'h0;
    font[815] = 8'h0;
    font[816] = 8'h0;
    font[817] = 8'h0;
    font[818] = 8'h3c;
    font[819] = 8'h42;
    font[820] = 8'h42;
    font[821] = 8'h2;
    font[822] = 8'h1c;
    font[823] = 8'h2;
    font[824] = 8'h2;
    font[825] = 8'h42;
    font[826] = 8'h42;
    font[827] = 8'h3c;
    font[828] = 8'h0;
    font[829] = 8'h0;
    font[830] = 8'h0;
    font[831] = 8'h0;
    font[832] = 8'h0;
    font[833] = 8'h0;
    font[834] = 8'h2;
    font[835] = 8'h6;
    font[836] = 8'ha;
    font[837] = 8'h12;
    font[838] = 8'h22;
    font[839] = 8'h42;
    font[840] = 8'h7e;
    font[841] = 8'h2;
    font[842] = 8'h2;
    font[843] = 8'h2;
    font[844] = 8'h0;
    font[845] = 8'h0;
    font[846] = 8'h0;
    font[847] = 8'h0;
    font[848] = 8'h0;
    font[849] = 8'h0;
    font[850] = 8'h7e;
    font[851] = 8'h40;
    font[852] = 8'h40;
    font[853] = 8'h40;
    font[854] = 8'h7c;
    font[855] = 8'h2;
    font[856] = 8'h2;
    font[857] = 8'h2;
    font[858] = 8'h42;
    font[859] = 8'h3c;
    font[860] = 8'h0;
    font[861] = 8'h0;
    font[862] = 8'h0;
    font[863] = 8'h0;
    font[864] = 8'h0;
    font[865] = 8'h0;
    font[866] = 8'h1c;
    font[867] = 8'h20;
    font[868] = 8'h40;
    font[869] = 8'h40;
    font[870] = 8'h7c;
    font[871] = 8'h42;
    font[872] = 8'h42;
    font[873] = 8'h42;
    font[874] = 8'h42;
    font[875] = 8'h3c;
    font[876] = 8'h0;
    font[877] = 8'h0;
    font[878] = 8'h0;
    font[879] = 8'h0;
    font[880] = 8'h0;
    font[881] = 8'h0;
    font[882] = 8'h7e;
    font[883] = 8'h2;
    font[884] = 8'h2;
    font[885] = 8'h4;
    font[886] = 8'h4;
    font[887] = 8'h8;
    font[888] = 8'h8;
    font[889] = 8'h10;
    font[890] = 8'h10;
    font[891] = 8'h10;
    font[892] = 8'h0;
    font[893] = 8'h0;
    font[894] = 8'h0;
    font[895] = 8'h0;
    font[896] = 8'h0;
    font[897] = 8'h0;
    font[898] = 8'h3c;
    font[899] = 8'h42;
    font[900] = 8'h42;
    font[901] = 8'h42;
    font[902] = 8'h3c;
    font[903] = 8'h42;
    font[904] = 8'h42;
    font[905] = 8'h42;
    font[906] = 8'h42;
    font[907] = 8'h3c;
    font[908] = 8'h0;
    font[909] = 8'h0;
    font[910] = 8'h0;
    font[911] = 8'h0;
    font[912] = 8'h0;
    font[913] = 8'h0;
    font[914] = 8'h3c;
    font[915] = 8'h42;
    font[916] = 8'h42;
    font[917] = 8'h42;
    font[918] = 8'h42;
    font[919] = 8'h3e;
    font[920] = 8'h2;
    font[921] = 8'h2;
    font[922] = 8'h4;
    font[923] = 8'h38;
    font[924] = 8'h0;
    font[925] = 8'h0;
    font[926] = 8'h0;
    font[927] = 8'h0;
    font[928] = 8'h0;
    font[929] = 8'h0;
    font[930] = 8'h0;
    font[931] = 8'h0;
    font[932] = 8'h0;
    font[933] = 8'h10;
    font[934] = 8'h10;
    font[935] = 8'h0;
    font[936] = 8'h0;
    font[937] = 8'h0;
    font[938] = 8'h10;
    font[939] = 8'h10;
    font[940] = 8'h0;
    font[941] = 8'h0;
    font[942] = 8'h0;
    font[943] = 8'h0;
    font[944] = 8'h0;
    font[945] = 8'h0;
    font[946] = 8'h0;
    font[947] = 8'h0;
    font[948] = 8'h0;
    font[949] = 8'h10;
    font[950] = 8'h10;
    font[951] = 8'h0;
    font[952] = 8'h0;
    font[953] = 8'h0;
    font[954] = 8'h10;
    font[955] = 8'h10;
    font[956] = 8'h20;
    font[957] = 8'h0;
    font[958] = 8'h0;
    font[959] = 8'h0;
    font[960] = 8'h0;
    font[961] = 8'h0;
    font[962] = 8'h0;
    font[963] = 8'h4;
    font[964] = 8'h8;
    font[965] = 8'h10;
    font[966] = 8'h20;
    font[967] = 8'h40;
    font[968] = 8'h20;
    font[969] = 8'h10;
    font[970] = 8'h8;
    font[971] = 8'h4;
    font[972] = 8'h0;
    font[973] = 8'h0;
    font[974] = 8'h0;
    font[975] = 8'h0;
    font[976] = 8'h0;
    font[977] = 8'h0;
    font[978] = 8'h0;
    font[979] = 8'h0;
    font[980] = 8'h0;
    font[981] = 8'h7e;
    font[982] = 8'h0;
    font[983] = 8'h0;
    font[984] = 8'h7e;
    font[985] = 8'h0;
    font[986] = 8'h0;
    font[987] = 8'h0;
    font[988] = 8'h0;
    font[989] = 8'h0;
    font[990] = 8'h0;
    font[991] = 8'h0;
    font[992] = 8'h0;
    font[993] = 8'h0;
    font[994] = 8'h0;
    font[995] = 8'h40;
    font[996] = 8'h20;
    font[997] = 8'h10;
    font[998] = 8'h8;
    font[999] = 8'h4;
    font[1000] = 8'h8;
    font[1001] = 8'h10;
    font[1002] = 8'h20;
    font[1003] = 8'h40;
    font[1004] = 8'h0;
    font[1005] = 8'h0;
    font[1006] = 8'h0;
    font[1007] = 8'h0;
    font[1008] = 8'h0;
    font[1009] = 8'h0;
    font[1010] = 8'h3c;
    font[1011] = 8'h42;
    font[1012] = 8'h42;
    font[1013] = 8'h42;
    font[1014] = 8'h4;
    font[1015] = 8'h8;
    font[1016] = 8'h8;
    font[1017] = 8'h0;
    font[1018] = 8'h8;
    font[1019] = 8'h8;
    font[1020] = 8'h0;
    font[1021] = 8'h0;
    font[1022] = 8'h0;
    font[1023] = 8'h0;
    font[1024] = 8'h0;
    font[1025] = 8'h0;
    font[1026] = 8'h7c;
    font[1027] = 8'h82;
    font[1028] = 8'h9e;
    font[1029] = 8'ha2;
    font[1030] = 8'ha2;
    font[1031] = 8'ha2;
    font[1032] = 8'ha6;
    font[1033] = 8'h9a;
    font[1034] = 8'h80;
    font[1035] = 8'h7e;
    font[1036] = 8'h0;
    font[1037] = 8'h0;
    font[1038] = 8'h0;
    font[1039] = 8'h0;
    font[1040] = 8'h0;
    font[1041] = 8'h0;
    font[1042] = 8'h3c;
    font[1043] = 8'h42;
    font[1044] = 8'h42;
    font[1045] = 8'h42;
    font[1046] = 8'h42;
    font[1047] = 8'h7e;
    font[1048] = 8'h42;
    font[1049] = 8'h42;
    font[1050] = 8'h42;
    font[1051] = 8'h42;
    font[1052] = 8'h0;
    font[1053] = 8'h0;
    font[1054] = 8'h0;
    font[1055] = 8'h0;
    font[1056] = 8'h0;
    font[1057] = 8'h0;
    font[1058] = 8'h7c;
    font[1059] = 8'h42;
    font[1060] = 8'h42;
    font[1061] = 8'h42;
    font[1062] = 8'h7c;
    font[1063] = 8'h42;
    font[1064] = 8'h42;
    font[1065] = 8'h42;
    font[1066] = 8'h42;
    font[1067] = 8'h7c;
    font[1068] = 8'h0;
    font[1069] = 8'h0;
    font[1070] = 8'h0;
    font[1071] = 8'h0;
    font[1072] = 8'h0;
    font[1073] = 8'h0;
    font[1074] = 8'h3c;
    font[1075] = 8'h42;
    font[1076] = 8'h42;
    font[1077] = 8'h40;
    font[1078] = 8'h40;
    font[1079] = 8'h40;
    font[1080] = 8'h40;
    font[1081] = 8'h42;
    font[1082] = 8'h42;
    font[1083] = 8'h3c;
    font[1084] = 8'h0;
    font[1085] = 8'h0;
    font[1086] = 8'h0;
    font[1087] = 8'h0;
    font[1088] = 8'h0;
    font[1089] = 8'h0;
    font[1090] = 8'h78;
    font[1091] = 8'h44;
    font[1092] = 8'h42;
    font[1093] = 8'h42;
    font[1094] = 8'h42;
    font[1095] = 8'h42;
    font[1096] = 8'h42;
    font[1097] = 8'h42;
    font[1098] = 8'h44;
    font[1099] = 8'h78;
    font[1100] = 8'h0;
    font[1101] = 8'h0;
    font[1102] = 8'h0;
    font[1103] = 8'h0;
    font[1104] = 8'h0;
    font[1105] = 8'h0;
    font[1106] = 8'h7e;
    font[1107] = 8'h40;
    font[1108] = 8'h40;
    font[1109] = 8'h40;
    font[1110] = 8'h78;
    font[1111] = 8'h40;
    font[1112] = 8'h40;
    font[1113] = 8'h40;
    font[1114] = 8'h40;
    font[1115] = 8'h7e;
    font[1116] = 8'h0;
    font[1117] = 8'h0;
    font[1118] = 8'h0;
    font[1119] = 8'h0;
    font[1120] = 8'h0;
    font[1121] = 8'h0;
    font[1122] = 8'h7e;
    font[1123] = 8'h40;
    font[1124] = 8'h40;
    font[1125] = 8'h40;
    font[1126] = 8'h78;
    font[1127] = 8'h40;
    font[1128] = 8'h40;
    font[1129] = 8'h40;
    font[1130] = 8'h40;
    font[1131] = 8'h40;
    font[1132] = 8'h0;
    font[1133] = 8'h0;
    font[1134] = 8'h0;
    font[1135] = 8'h0;
    font[1136] = 8'h0;
    font[1137] = 8'h0;
    font[1138] = 8'h3c;
    font[1139] = 8'h42;
    font[1140] = 8'h42;
    font[1141] = 8'h40;
    font[1142] = 8'h40;
    font[1143] = 8'h4e;
    font[1144] = 8'h42;
    font[1145] = 8'h42;
    font[1146] = 8'h42;
    font[1147] = 8'h3c;
    font[1148] = 8'h0;
    font[1149] = 8'h0;
    font[1150] = 8'h0;
    font[1151] = 8'h0;
    font[1152] = 8'h0;
    font[1153] = 8'h0;
    font[1154] = 8'h42;
    font[1155] = 8'h42;
    font[1156] = 8'h42;
    font[1157] = 8'h42;
    font[1158] = 8'h7e;
    font[1159] = 8'h42;
    font[1160] = 8'h42;
    font[1161] = 8'h42;
    font[1162] = 8'h42;
    font[1163] = 8'h42;
    font[1164] = 8'h0;
    font[1165] = 8'h0;
    font[1166] = 8'h0;
    font[1167] = 8'h0;
    font[1168] = 8'h0;
    font[1169] = 8'h0;
    font[1170] = 8'h38;
    font[1171] = 8'h10;
    font[1172] = 8'h10;
    font[1173] = 8'h10;
    font[1174] = 8'h10;
    font[1175] = 8'h10;
    font[1176] = 8'h10;
    font[1177] = 8'h10;
    font[1178] = 8'h10;
    font[1179] = 8'h38;
    font[1180] = 8'h0;
    font[1181] = 8'h0;
    font[1182] = 8'h0;
    font[1183] = 8'h0;
    font[1184] = 8'h0;
    font[1185] = 8'h0;
    font[1186] = 8'he;
    font[1187] = 8'h4;
    font[1188] = 8'h4;
    font[1189] = 8'h4;
    font[1190] = 8'h4;
    font[1191] = 8'h4;
    font[1192] = 8'h4;
    font[1193] = 8'h44;
    font[1194] = 8'h44;
    font[1195] = 8'h38;
    font[1196] = 8'h0;
    font[1197] = 8'h0;
    font[1198] = 8'h0;
    font[1199] = 8'h0;
    font[1200] = 8'h0;
    font[1201] = 8'h0;
    font[1202] = 8'h42;
    font[1203] = 8'h44;
    font[1204] = 8'h48;
    font[1205] = 8'h50;
    font[1206] = 8'h60;
    font[1207] = 8'h60;
    font[1208] = 8'h50;
    font[1209] = 8'h48;
    font[1210] = 8'h44;
    font[1211] = 8'h42;
    font[1212] = 8'h0;
    font[1213] = 8'h0;
    font[1214] = 8'h0;
    font[1215] = 8'h0;
    font[1216] = 8'h0;
    font[1217] = 8'h0;
    font[1218] = 8'h40;
    font[1219] = 8'h40;
    font[1220] = 8'h40;
    font[1221] = 8'h40;
    font[1222] = 8'h40;
    font[1223] = 8'h40;
    font[1224] = 8'h40;
    font[1225] = 8'h40;
    font[1226] = 8'h40;
    font[1227] = 8'h7e;
    font[1228] = 8'h0;
    font[1229] = 8'h0;
    font[1230] = 8'h0;
    font[1231] = 8'h0;
    font[1232] = 8'h0;
    font[1233] = 8'h0;
    font[1234] = 8'h82;
    font[1235] = 8'hc6;
    font[1236] = 8'haa;
    font[1237] = 8'h92;
    font[1238] = 8'h92;
    font[1239] = 8'h82;
    font[1240] = 8'h82;
    font[1241] = 8'h82;
    font[1242] = 8'h82;
    font[1243] = 8'h82;
    font[1244] = 8'h0;
    font[1245] = 8'h0;
    font[1246] = 8'h0;
    font[1247] = 8'h0;
    font[1248] = 8'h0;
    font[1249] = 8'h0;
    font[1250] = 8'h42;
    font[1251] = 8'h42;
    font[1252] = 8'h42;
    font[1253] = 8'h62;
    font[1254] = 8'h52;
    font[1255] = 8'h4a;
    font[1256] = 8'h46;
    font[1257] = 8'h42;
    font[1258] = 8'h42;
    font[1259] = 8'h42;
    font[1260] = 8'h0;
    font[1261] = 8'h0;
    font[1262] = 8'h0;
    font[1263] = 8'h0;
    font[1264] = 8'h0;
    font[1265] = 8'h0;
    font[1266] = 8'h3c;
    font[1267] = 8'h42;
    font[1268] = 8'h42;
    font[1269] = 8'h42;
    font[1270] = 8'h42;
    font[1271] = 8'h42;
    font[1272] = 8'h42;
    font[1273] = 8'h42;
    font[1274] = 8'h42;
    font[1275] = 8'h3c;
    font[1276] = 8'h0;
    font[1277] = 8'h0;
    font[1278] = 8'h0;
    font[1279] = 8'h0;
    font[1280] = 8'h0;
    font[1281] = 8'h0;
    font[1282] = 8'h7c;
    font[1283] = 8'h42;
    font[1284] = 8'h42;
    font[1285] = 8'h42;
    font[1286] = 8'h42;
    font[1287] = 8'h7c;
    font[1288] = 8'h40;
    font[1289] = 8'h40;
    font[1290] = 8'h40;
    font[1291] = 8'h40;
    font[1292] = 8'h0;
    font[1293] = 8'h0;
    font[1294] = 8'h0;
    font[1295] = 8'h0;
    font[1296] = 8'h0;
    font[1297] = 8'h0;
    font[1298] = 8'h3c;
    font[1299] = 8'h42;
    font[1300] = 8'h42;
    font[1301] = 8'h42;
    font[1302] = 8'h42;
    font[1303] = 8'h42;
    font[1304] = 8'h42;
    font[1305] = 8'h42;
    font[1306] = 8'h4a;
    font[1307] = 8'h3c;
    font[1308] = 8'h2;
    font[1309] = 8'h0;
    font[1310] = 8'h0;
    font[1311] = 8'h0;
    font[1312] = 8'h0;
    font[1313] = 8'h0;
    font[1314] = 8'h7c;
    font[1315] = 8'h42;
    font[1316] = 8'h42;
    font[1317] = 8'h42;
    font[1318] = 8'h42;
    font[1319] = 8'h7c;
    font[1320] = 8'h50;
    font[1321] = 8'h48;
    font[1322] = 8'h44;
    font[1323] = 8'h42;
    font[1324] = 8'h0;
    font[1325] = 8'h0;
    font[1326] = 8'h0;
    font[1327] = 8'h0;
    font[1328] = 8'h0;
    font[1329] = 8'h0;
    font[1330] = 8'h3c;
    font[1331] = 8'h42;
    font[1332] = 8'h40;
    font[1333] = 8'h40;
    font[1334] = 8'h3c;
    font[1335] = 8'h2;
    font[1336] = 8'h2;
    font[1337] = 8'h42;
    font[1338] = 8'h42;
    font[1339] = 8'h3c;
    font[1340] = 8'h0;
    font[1341] = 8'h0;
    font[1342] = 8'h0;
    font[1343] = 8'h0;
    font[1344] = 8'h0;
    font[1345] = 8'h0;
    font[1346] = 8'hfe;
    font[1347] = 8'h10;
    font[1348] = 8'h10;
    font[1349] = 8'h10;
    font[1350] = 8'h10;
    font[1351] = 8'h10;
    font[1352] = 8'h10;
    font[1353] = 8'h10;
    font[1354] = 8'h10;
    font[1355] = 8'h10;
    font[1356] = 8'h0;
    font[1357] = 8'h0;
    font[1358] = 8'h0;
    font[1359] = 8'h0;
    font[1360] = 8'h0;
    font[1361] = 8'h0;
    font[1362] = 8'h42;
    font[1363] = 8'h42;
    font[1364] = 8'h42;
    font[1365] = 8'h42;
    font[1366] = 8'h42;
    font[1367] = 8'h42;
    font[1368] = 8'h42;
    font[1369] = 8'h42;
    font[1370] = 8'h42;
    font[1371] = 8'h3c;
    font[1372] = 8'h0;
    font[1373] = 8'h0;
    font[1374] = 8'h0;
    font[1375] = 8'h0;
    font[1376] = 8'h0;
    font[1377] = 8'h0;
    font[1378] = 8'h42;
    font[1379] = 8'h42;
    font[1380] = 8'h42;
    font[1381] = 8'h42;
    font[1382] = 8'h42;
    font[1383] = 8'h24;
    font[1384] = 8'h24;
    font[1385] = 8'h24;
    font[1386] = 8'h18;
    font[1387] = 8'h18;
    font[1388] = 8'h0;
    font[1389] = 8'h0;
    font[1390] = 8'h0;
    font[1391] = 8'h0;
    font[1392] = 8'h0;
    font[1393] = 8'h0;
    font[1394] = 8'h82;
    font[1395] = 8'h82;
    font[1396] = 8'h82;
    font[1397] = 8'h82;
    font[1398] = 8'h82;
    font[1399] = 8'h92;
    font[1400] = 8'h92;
    font[1401] = 8'haa;
    font[1402] = 8'hc6;
    font[1403] = 8'h82;
    font[1404] = 8'h0;
    font[1405] = 8'h0;
    font[1406] = 8'h0;
    font[1407] = 8'h0;
    font[1408] = 8'h0;
    font[1409] = 8'h0;
    font[1410] = 8'h42;
    font[1411] = 8'h42;
    font[1412] = 8'h24;
    font[1413] = 8'h24;
    font[1414] = 8'h18;
    font[1415] = 8'h18;
    font[1416] = 8'h24;
    font[1417] = 8'h24;
    font[1418] = 8'h42;
    font[1419] = 8'h42;
    font[1420] = 8'h0;
    font[1421] = 8'h0;
    font[1422] = 8'h0;
    font[1423] = 8'h0;
    font[1424] = 8'h0;
    font[1425] = 8'h0;
    font[1426] = 8'h82;
    font[1427] = 8'h82;
    font[1428] = 8'h44;
    font[1429] = 8'h44;
    font[1430] = 8'h28;
    font[1431] = 8'h10;
    font[1432] = 8'h10;
    font[1433] = 8'h10;
    font[1434] = 8'h10;
    font[1435] = 8'h10;
    font[1436] = 8'h0;
    font[1437] = 8'h0;
    font[1438] = 8'h0;
    font[1439] = 8'h0;
    font[1440] = 8'h0;
    font[1441] = 8'h0;
    font[1442] = 8'h7e;
    font[1443] = 8'h2;
    font[1444] = 8'h2;
    font[1445] = 8'h4;
    font[1446] = 8'h8;
    font[1447] = 8'h10;
    font[1448] = 8'h20;
    font[1449] = 8'h40;
    font[1450] = 8'h40;
    font[1451] = 8'h7e;
    font[1452] = 8'h0;
    font[1453] = 8'h0;
    font[1454] = 8'h0;
    font[1455] = 8'h0;
    font[1456] = 8'h0;
    font[1457] = 8'h0;
    font[1458] = 8'h38;
    font[1459] = 8'h20;
    font[1460] = 8'h20;
    font[1461] = 8'h20;
    font[1462] = 8'h20;
    font[1463] = 8'h20;
    font[1464] = 8'h20;
    font[1465] = 8'h20;
    font[1466] = 8'h20;
    font[1467] = 8'h38;
    font[1468] = 8'h0;
    font[1469] = 8'h0;
    font[1470] = 8'h0;
    font[1471] = 8'h0;
    font[1472] = 8'h0;
    font[1473] = 8'h0;
    font[1474] = 8'h40;
    font[1475] = 8'h40;
    font[1476] = 8'h20;
    font[1477] = 8'h20;
    font[1478] = 8'h10;
    font[1479] = 8'h10;
    font[1480] = 8'h8;
    font[1481] = 8'h8;
    font[1482] = 8'h4;
    font[1483] = 8'h4;
    font[1484] = 8'h0;
    font[1485] = 8'h0;
    font[1486] = 8'h0;
    font[1487] = 8'h0;
    font[1488] = 8'h0;
    font[1489] = 8'h0;
    font[1490] = 8'h38;
    font[1491] = 8'h8;
    font[1492] = 8'h8;
    font[1493] = 8'h8;
    font[1494] = 8'h8;
    font[1495] = 8'h8;
    font[1496] = 8'h8;
    font[1497] = 8'h8;
    font[1498] = 8'h8;
    font[1499] = 8'h38;
    font[1500] = 8'h0;
    font[1501] = 8'h0;
    font[1502] = 8'h0;
    font[1503] = 8'h0;
    font[1504] = 8'h0;
    font[1505] = 8'h10;
    font[1506] = 8'h28;
    font[1507] = 8'h44;
    font[1508] = 8'h0;
    font[1509] = 8'h0;
    font[1510] = 8'h0;
    font[1511] = 8'h0;
    font[1512] = 8'h0;
    font[1513] = 8'h0;
    font[1514] = 8'h0;
    font[1515] = 8'h0;
    font[1516] = 8'h0;
    font[1517] = 8'h0;
    font[1518] = 8'h0;
    font[1519] = 8'h0;
    font[1520] = 8'h0;
    font[1521] = 8'h0;
    font[1522] = 8'h0;
    font[1523] = 8'h0;
    font[1524] = 8'h0;
    font[1525] = 8'h0;
    font[1526] = 8'h0;
    font[1527] = 8'h0;
    font[1528] = 8'h0;
    font[1529] = 8'h0;
    font[1530] = 8'h0;
    font[1531] = 8'h0;
    font[1532] = 8'h0;
    font[1533] = 8'h7e;
    font[1534] = 8'h0;
    font[1535] = 8'h0;
    font[1536] = 8'h10;
    font[1537] = 8'h8;
    font[1538] = 8'h0;
    font[1539] = 8'h0;
    font[1540] = 8'h0;
    font[1541] = 8'h0;
    font[1542] = 8'h0;
    font[1543] = 8'h0;
    font[1544] = 8'h0;
    font[1545] = 8'h0;
    font[1546] = 8'h0;
    font[1547] = 8'h0;
    font[1548] = 8'h0;
    font[1549] = 8'h0;
    font[1550] = 8'h0;
    font[1551] = 8'h0;
    font[1552] = 8'h0;
    font[1553] = 8'h0;
    font[1554] = 8'h0;
    font[1555] = 8'h0;
    font[1556] = 8'h0;
    font[1557] = 8'h3c;
    font[1558] = 8'h2;
    font[1559] = 8'h3e;
    font[1560] = 8'h42;
    font[1561] = 8'h42;
    font[1562] = 8'h42;
    font[1563] = 8'h3e;
    font[1564] = 8'h0;
    font[1565] = 8'h0;
    font[1566] = 8'h0;
    font[1567] = 8'h0;
    font[1568] = 8'h0;
    font[1569] = 8'h0;
    font[1570] = 8'h40;
    font[1571] = 8'h40;
    font[1572] = 8'h40;
    font[1573] = 8'h7c;
    font[1574] = 8'h42;
    font[1575] = 8'h42;
    font[1576] = 8'h42;
    font[1577] = 8'h42;
    font[1578] = 8'h42;
    font[1579] = 8'h7c;
    font[1580] = 8'h0;
    font[1581] = 8'h0;
    font[1582] = 8'h0;
    font[1583] = 8'h0;
    font[1584] = 8'h0;
    font[1585] = 8'h0;
    font[1586] = 8'h0;
    font[1587] = 8'h0;
    font[1588] = 8'h0;
    font[1589] = 8'h3c;
    font[1590] = 8'h42;
    font[1591] = 8'h40;
    font[1592] = 8'h40;
    font[1593] = 8'h40;
    font[1594] = 8'h42;
    font[1595] = 8'h3c;
    font[1596] = 8'h0;
    font[1597] = 8'h0;
    font[1598] = 8'h0;
    font[1599] = 8'h0;
    font[1600] = 8'h0;
    font[1601] = 8'h0;
    font[1602] = 8'h2;
    font[1603] = 8'h2;
    font[1604] = 8'h2;
    font[1605] = 8'h3e;
    font[1606] = 8'h42;
    font[1607] = 8'h42;
    font[1608] = 8'h42;
    font[1609] = 8'h42;
    font[1610] = 8'h42;
    font[1611] = 8'h3e;
    font[1612] = 8'h0;
    font[1613] = 8'h0;
    font[1614] = 8'h0;
    font[1615] = 8'h0;
    font[1616] = 8'h0;
    font[1617] = 8'h0;
    font[1618] = 8'h0;
    font[1619] = 8'h0;
    font[1620] = 8'h0;
    font[1621] = 8'h3c;
    font[1622] = 8'h42;
    font[1623] = 8'h42;
    font[1624] = 8'h7e;
    font[1625] = 8'h40;
    font[1626] = 8'h40;
    font[1627] = 8'h3c;
    font[1628] = 8'h0;
    font[1629] = 8'h0;
    font[1630] = 8'h0;
    font[1631] = 8'h0;
    font[1632] = 8'h0;
    font[1633] = 8'h0;
    font[1634] = 8'he;
    font[1635] = 8'h10;
    font[1636] = 8'h10;
    font[1637] = 8'h7c;
    font[1638] = 8'h10;
    font[1639] = 8'h10;
    font[1640] = 8'h10;
    font[1641] = 8'h10;
    font[1642] = 8'h10;
    font[1643] = 8'h10;
    font[1644] = 8'h0;
    font[1645] = 8'h0;
    font[1646] = 8'h0;
    font[1647] = 8'h0;
    font[1648] = 8'h0;
    font[1649] = 8'h0;
    font[1650] = 8'h0;
    font[1651] = 8'h0;
    font[1652] = 8'h0;
    font[1653] = 8'h3e;
    font[1654] = 8'h42;
    font[1655] = 8'h42;
    font[1656] = 8'h42;
    font[1657] = 8'h42;
    font[1658] = 8'h42;
    font[1659] = 8'h3e;
    font[1660] = 8'h2;
    font[1661] = 8'h2;
    font[1662] = 8'h3c;
    font[1663] = 8'h0;
    font[1664] = 8'h0;
    font[1665] = 8'h0;
    font[1666] = 8'h40;
    font[1667] = 8'h40;
    font[1668] = 8'h40;
    font[1669] = 8'h7c;
    font[1670] = 8'h42;
    font[1671] = 8'h42;
    font[1672] = 8'h42;
    font[1673] = 8'h42;
    font[1674] = 8'h42;
    font[1675] = 8'h42;
    font[1676] = 8'h0;
    font[1677] = 8'h0;
    font[1678] = 8'h0;
    font[1679] = 8'h0;
    font[1680] = 8'h0;
    font[1681] = 8'h0;
    font[1682] = 8'h10;
    font[1683] = 8'h10;
    font[1684] = 8'h0;
    font[1685] = 8'h30;
    font[1686] = 8'h10;
    font[1687] = 8'h10;
    font[1688] = 8'h10;
    font[1689] = 8'h10;
    font[1690] = 8'h10;
    font[1691] = 8'h38;
    font[1692] = 8'h0;
    font[1693] = 8'h0;
    font[1694] = 8'h0;
    font[1695] = 8'h0;
    font[1696] = 8'h0;
    font[1697] = 8'h0;
    font[1698] = 8'h4;
    font[1699] = 8'h4;
    font[1700] = 8'h0;
    font[1701] = 8'hc;
    font[1702] = 8'h4;
    font[1703] = 8'h4;
    font[1704] = 8'h4;
    font[1705] = 8'h4;
    font[1706] = 8'h4;
    font[1707] = 8'h4;
    font[1708] = 8'h44;
    font[1709] = 8'h44;
    font[1710] = 8'h38;
    font[1711] = 8'h0;
    font[1712] = 8'h0;
    font[1713] = 8'h0;
    font[1714] = 8'h40;
    font[1715] = 8'h40;
    font[1716] = 8'h40;
    font[1717] = 8'h42;
    font[1718] = 8'h44;
    font[1719] = 8'h48;
    font[1720] = 8'h70;
    font[1721] = 8'h48;
    font[1722] = 8'h44;
    font[1723] = 8'h42;
    font[1724] = 8'h0;
    font[1725] = 8'h0;
    font[1726] = 8'h0;
    font[1727] = 8'h0;
    font[1728] = 8'h0;
    font[1729] = 8'h0;
    font[1730] = 8'h30;
    font[1731] = 8'h10;
    font[1732] = 8'h10;
    font[1733] = 8'h10;
    font[1734] = 8'h10;
    font[1735] = 8'h10;
    font[1736] = 8'h10;
    font[1737] = 8'h10;
    font[1738] = 8'h10;
    font[1739] = 8'h38;
    font[1740] = 8'h0;
    font[1741] = 8'h0;
    font[1742] = 8'h0;
    font[1743] = 8'h0;
    font[1744] = 8'h0;
    font[1745] = 8'h0;
    font[1746] = 8'h0;
    font[1747] = 8'h0;
    font[1748] = 8'h0;
    font[1749] = 8'hfc;
    font[1750] = 8'h92;
    font[1751] = 8'h92;
    font[1752] = 8'h92;
    font[1753] = 8'h92;
    font[1754] = 8'h92;
    font[1755] = 8'h92;
    font[1756] = 8'h0;
    font[1757] = 8'h0;
    font[1758] = 8'h0;
    font[1759] = 8'h0;
    font[1760] = 8'h0;
    font[1761] = 8'h0;
    font[1762] = 8'h0;
    font[1763] = 8'h0;
    font[1764] = 8'h0;
    font[1765] = 8'h7c;
    font[1766] = 8'h42;
    font[1767] = 8'h42;
    font[1768] = 8'h42;
    font[1769] = 8'h42;
    font[1770] = 8'h42;
    font[1771] = 8'h42;
    font[1772] = 8'h0;
    font[1773] = 8'h0;
    font[1774] = 8'h0;
    font[1775] = 8'h0;
    font[1776] = 8'h0;
    font[1777] = 8'h0;
    font[1778] = 8'h0;
    font[1779] = 8'h0;
    font[1780] = 8'h0;
    font[1781] = 8'h3c;
    font[1782] = 8'h42;
    font[1783] = 8'h42;
    font[1784] = 8'h42;
    font[1785] = 8'h42;
    font[1786] = 8'h42;
    font[1787] = 8'h3c;
    font[1788] = 8'h0;
    font[1789] = 8'h0;
    font[1790] = 8'h0;
    font[1791] = 8'h0;
    font[1792] = 8'h0;
    font[1793] = 8'h0;
    font[1794] = 8'h0;
    font[1795] = 8'h0;
    font[1796] = 8'h0;
    font[1797] = 8'h7c;
    font[1798] = 8'h42;
    font[1799] = 8'h42;
    font[1800] = 8'h42;
    font[1801] = 8'h42;
    font[1802] = 8'h42;
    font[1803] = 8'h7c;
    font[1804] = 8'h40;
    font[1805] = 8'h40;
    font[1806] = 8'h40;
    font[1807] = 8'h0;
    font[1808] = 8'h0;
    font[1809] = 8'h0;
    font[1810] = 8'h0;
    font[1811] = 8'h0;
    font[1812] = 8'h0;
    font[1813] = 8'h3e;
    font[1814] = 8'h42;
    font[1815] = 8'h42;
    font[1816] = 8'h42;
    font[1817] = 8'h42;
    font[1818] = 8'h42;
    font[1819] = 8'h3e;
    font[1820] = 8'h2;
    font[1821] = 8'h2;
    font[1822] = 8'h2;
    font[1823] = 8'h0;
    font[1824] = 8'h0;
    font[1825] = 8'h0;
    font[1826] = 8'h0;
    font[1827] = 8'h0;
    font[1828] = 8'h0;
    font[1829] = 8'h5e;
    font[1830] = 8'h60;
    font[1831] = 8'h40;
    font[1832] = 8'h40;
    font[1833] = 8'h40;
    font[1834] = 8'h40;
    font[1835] = 8'h40;
    font[1836] = 8'h0;
    font[1837] = 8'h0;
    font[1838] = 8'h0;
    font[1839] = 8'h0;
    font[1840] = 8'h0;
    font[1841] = 8'h0;
    font[1842] = 8'h0;
    font[1843] = 8'h0;
    font[1844] = 8'h0;
    font[1845] = 8'h3e;
    font[1846] = 8'h40;
    font[1847] = 8'h40;
    font[1848] = 8'h3c;
    font[1849] = 8'h2;
    font[1850] = 8'h2;
    font[1851] = 8'h7c;
    font[1852] = 8'h0;
    font[1853] = 8'h0;
    font[1854] = 8'h0;
    font[1855] = 8'h0;
    font[1856] = 8'h0;
    font[1857] = 8'h0;
    font[1858] = 8'h10;
    font[1859] = 8'h10;
    font[1860] = 8'h10;
    font[1861] = 8'h7c;
    font[1862] = 8'h10;
    font[1863] = 8'h10;
    font[1864] = 8'h10;
    font[1865] = 8'h10;
    font[1866] = 8'h10;
    font[1867] = 8'he;
    font[1868] = 8'h0;
    font[1869] = 8'h0;
    font[1870] = 8'h0;
    font[1871] = 8'h0;
    font[1872] = 8'h0;
    font[1873] = 8'h0;
    font[1874] = 8'h0;
    font[1875] = 8'h0;
    font[1876] = 8'h0;
    font[1877] = 8'h42;
    font[1878] = 8'h42;
    font[1879] = 8'h42;
    font[1880] = 8'h42;
    font[1881] = 8'h42;
    font[1882] = 8'h42;
    font[1883] = 8'h3e;
    font[1884] = 8'h0;
    font[1885] = 8'h0;
    font[1886] = 8'h0;
    font[1887] = 8'h0;
    font[1888] = 8'h0;
    font[1889] = 8'h0;
    font[1890] = 8'h0;
    font[1891] = 8'h0;
    font[1892] = 8'h0;
    font[1893] = 8'h42;
    font[1894] = 8'h42;
    font[1895] = 8'h42;
    font[1896] = 8'h24;
    font[1897] = 8'h24;
    font[1898] = 8'h18;
    font[1899] = 8'h18;
    font[1900] = 8'h0;
    font[1901] = 8'h0;
    font[1902] = 8'h0;
    font[1903] = 8'h0;
    font[1904] = 8'h0;
    font[1905] = 8'h0;
    font[1906] = 8'h0;
    font[1907] = 8'h0;
    font[1908] = 8'h0;
    font[1909] = 8'h82;
    font[1910] = 8'h82;
    font[1911] = 8'h92;
    font[1912] = 8'h92;
    font[1913] = 8'h92;
    font[1914] = 8'h92;
    font[1915] = 8'h7c;
    font[1916] = 8'h0;
    font[1917] = 8'h0;
    font[1918] = 8'h0;
    font[1919] = 8'h0;
    font[1920] = 8'h0;
    font[1921] = 8'h0;
    font[1922] = 8'h0;
    font[1923] = 8'h0;
    font[1924] = 8'h0;
    font[1925] = 8'h42;
    font[1926] = 8'h42;
    font[1927] = 8'h24;
    font[1928] = 8'h18;
    font[1929] = 8'h24;
    font[1930] = 8'h42;
    font[1931] = 8'h42;
    font[1932] = 8'h0;
    font[1933] = 8'h0;
    font[1934] = 8'h0;
    font[1935] = 8'h0;
    font[1936] = 8'h0;
    font[1937] = 8'h0;
    font[1938] = 8'h0;
    font[1939] = 8'h0;
    font[1940] = 8'h0;
    font[1941] = 8'h42;
    font[1942] = 8'h42;
    font[1943] = 8'h42;
    font[1944] = 8'h42;
    font[1945] = 8'h42;
    font[1946] = 8'h42;
    font[1947] = 8'h3e;
    font[1948] = 8'h2;
    font[1949] = 8'h2;
    font[1950] = 8'h3c;
    font[1951] = 8'h0;
    font[1952] = 8'h0;
    font[1953] = 8'h0;
    font[1954] = 8'h0;
    font[1955] = 8'h0;
    font[1956] = 8'h0;
    font[1957] = 8'h7e;
    font[1958] = 8'h4;
    font[1959] = 8'h8;
    font[1960] = 8'h10;
    font[1961] = 8'h20;
    font[1962] = 8'h40;
    font[1963] = 8'h7e;
    font[1964] = 8'h0;
    font[1965] = 8'h0;
    font[1966] = 8'h0;
    font[1967] = 8'h0;
    font[1968] = 8'h0;
    font[1969] = 8'h0;
    font[1970] = 8'hc;
    font[1971] = 8'h10;
    font[1972] = 8'h10;
    font[1973] = 8'h10;
    font[1974] = 8'h20;
    font[1975] = 8'h10;
    font[1976] = 8'h10;
    font[1977] = 8'h10;
    font[1978] = 8'h10;
    font[1979] = 8'hc;
    font[1980] = 8'h0;
    font[1981] = 8'h0;
    font[1982] = 8'h0;
    font[1983] = 8'h0;
    font[1984] = 8'h0;
    font[1985] = 8'h0;
    font[1986] = 8'h10;
    font[1987] = 8'h10;
    font[1988] = 8'h10;
    font[1989] = 8'h10;
    font[1990] = 8'h10;
    font[1991] = 8'h10;
    font[1992] = 8'h10;
    font[1993] = 8'h10;
    font[1994] = 8'h10;
    font[1995] = 8'h10;
    font[1996] = 8'h0;
    font[1997] = 8'h0;
    font[1998] = 8'h0;
    font[1999] = 8'h0;
    font[2000] = 8'h0;
    font[2001] = 8'h0;
    font[2002] = 8'h30;
    font[2003] = 8'h8;
    font[2004] = 8'h8;
    font[2005] = 8'h8;
    font[2006] = 8'h4;
    font[2007] = 8'h8;
    font[2008] = 8'h8;
    font[2009] = 8'h8;
    font[2010] = 8'h8;
    font[2011] = 8'h30;
    font[2012] = 8'h0;
    font[2013] = 8'h0;
    font[2014] = 8'h0;
    font[2015] = 8'h0;
    font[2016] = 8'h0;
    font[2017] = 8'h62;
    font[2018] = 8'h92;
    font[2019] = 8'h8c;
  end
endmodule
